// Dummy implementation, does nothing
module TC_SegmentDisplay (clk, rst, enable, value);
    parameter UUID = 0;
    parameter NAME = "";
    input clk;
    input rst;
    input enable;
    input [7:0] value;
endmodule
