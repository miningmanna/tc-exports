
module TC_Clock(clk, rst);
    parameter UUID = 0;
    parameter NAME = "";
    output out;
    
    assign out = clk;
endmodule
